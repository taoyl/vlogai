interface example_mod (
    axi4mst cpucore_mst
   ,axi4slv syscsr_slv
   ,.*
);
endinterface
